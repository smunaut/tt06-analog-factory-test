magic
tech sky130A
magscale 1 2
timestamp 1713640305
<< locali >>
rect 5024 38334 11630 38410
rect 5024 38286 5036 38334
rect 11618 38286 11630 38334
rect 5024 38280 11630 38286
<< viali >>
rect 5036 38286 11618 38334
<< metal1 >>
rect 11070 39146 11136 39152
rect 5040 39140 5108 39146
rect 5040 39086 5046 39140
rect 5102 39086 5108 39140
rect 5040 39080 5108 39086
rect 5518 39140 5584 39146
rect 5518 39086 5524 39140
rect 5578 39086 5584 39140
rect 11070 39092 11076 39146
rect 11130 39092 11136 39146
rect 11070 39086 11136 39092
rect 11544 39140 11612 39146
rect 11544 39086 11550 39140
rect 11606 39086 11612 39140
rect 5518 39080 5584 39086
rect 5056 39022 5090 39080
rect 5544 39022 5578 39080
rect 11076 39022 11110 39086
rect 11544 39080 11612 39086
rect 11560 39022 11594 39080
rect 5056 38988 5508 39022
rect 5056 38512 5090 38988
rect 5124 38936 5178 38950
rect 5124 38546 5178 38556
rect 5256 38944 5310 38950
rect 5256 38550 5310 38556
rect 5386 38936 5440 38950
rect 5386 38546 5440 38556
rect 5474 38512 5508 38988
rect 5056 38478 5508 38512
rect 5544 38988 11110 39022
rect 5544 38512 5578 38988
rect 5612 38940 5666 38950
rect 5612 38550 5666 38560
rect 5740 38940 5794 38950
rect 5740 38550 5794 38560
rect 5868 38940 5922 38950
rect 5868 38550 5922 38560
rect 5996 38940 6050 38950
rect 5996 38550 6050 38560
rect 6124 38940 6178 38950
rect 6124 38550 6178 38560
rect 6252 38940 6306 38950
rect 6252 38550 6306 38560
rect 6380 38940 6434 38950
rect 6380 38550 6434 38560
rect 6508 38940 6562 38950
rect 6508 38550 6562 38560
rect 6636 38940 6690 38950
rect 6636 38550 6690 38560
rect 6764 38940 6818 38950
rect 6764 38550 6818 38560
rect 6892 38940 6946 38950
rect 6892 38550 6946 38560
rect 7020 38940 7074 38950
rect 7020 38550 7074 38560
rect 7148 38940 7202 38950
rect 7148 38550 7202 38560
rect 7276 38940 7330 38950
rect 7276 38550 7330 38560
rect 7404 38940 7458 38950
rect 7404 38550 7458 38560
rect 7532 38940 7586 38950
rect 7532 38550 7586 38560
rect 7660 38940 7714 38950
rect 7660 38550 7714 38560
rect 7788 38940 7842 38950
rect 7788 38550 7842 38560
rect 7916 38940 7970 38950
rect 7916 38550 7970 38560
rect 8038 38512 8104 38988
rect 8172 38940 8226 38950
rect 8172 38550 8226 38560
rect 8300 38940 8354 38950
rect 8300 38550 8354 38560
rect 8428 38940 8482 38950
rect 8428 38550 8482 38560
rect 8556 38940 8610 38950
rect 8556 38550 8610 38560
rect 8684 38940 8738 38950
rect 8684 38550 8738 38560
rect 8812 38940 8866 38950
rect 8812 38550 8866 38560
rect 8940 38940 8994 38950
rect 8940 38550 8994 38560
rect 9068 38940 9122 38950
rect 9068 38550 9122 38560
rect 9196 38940 9250 38950
rect 9196 38550 9250 38560
rect 9324 38940 9378 38950
rect 9324 38550 9378 38560
rect 9452 38940 9506 38950
rect 9452 38550 9506 38560
rect 9580 38940 9634 38950
rect 9580 38550 9634 38560
rect 9708 38940 9762 38950
rect 9708 38550 9762 38560
rect 9836 38940 9890 38950
rect 9836 38550 9890 38560
rect 9964 38940 10018 38950
rect 9964 38550 10018 38560
rect 10092 38940 10146 38950
rect 10092 38550 10146 38560
rect 10220 38940 10274 38950
rect 10220 38550 10274 38560
rect 10348 38940 10402 38950
rect 10348 38550 10402 38560
rect 10476 38940 10530 38950
rect 10476 38550 10530 38560
rect 10604 38940 10658 38950
rect 10604 38550 10658 38560
rect 10732 38940 10786 38950
rect 10732 38550 10786 38560
rect 10860 38940 10914 38950
rect 10860 38550 10914 38560
rect 10988 38940 11042 38950
rect 10988 38550 11042 38560
rect 11076 38512 11110 38988
rect 5544 38478 11110 38512
rect 11148 38988 11594 39022
rect 11148 38512 11182 38988
rect 11216 38944 11270 38950
rect 11216 38550 11270 38556
rect 11344 38944 11398 38950
rect 11344 38550 11398 38556
rect 11472 38944 11526 38950
rect 11472 38550 11526 38556
rect 11560 38512 11594 38988
rect 11148 38478 11594 38512
rect 5024 38280 5030 38340
rect 11624 38280 11630 38340
<< via1 >>
rect 5046 39086 5102 39140
rect 5524 39086 5578 39140
rect 11076 39092 11130 39146
rect 11550 39086 11606 39140
rect 5124 38556 5178 38936
rect 5256 38556 5310 38944
rect 5386 38556 5440 38936
rect 5612 38560 5666 38940
rect 5740 38560 5794 38940
rect 5868 38560 5922 38940
rect 5996 38560 6050 38940
rect 6124 38560 6178 38940
rect 6252 38560 6306 38940
rect 6380 38560 6434 38940
rect 6508 38560 6562 38940
rect 6636 38560 6690 38940
rect 6764 38560 6818 38940
rect 6892 38560 6946 38940
rect 7020 38560 7074 38940
rect 7148 38560 7202 38940
rect 7276 38560 7330 38940
rect 7404 38560 7458 38940
rect 7532 38560 7586 38940
rect 7660 38560 7714 38940
rect 7788 38560 7842 38940
rect 7916 38560 7970 38940
rect 8172 38560 8226 38940
rect 8300 38560 8354 38940
rect 8428 38560 8482 38940
rect 8556 38560 8610 38940
rect 8684 38560 8738 38940
rect 8812 38560 8866 38940
rect 8940 38560 8994 38940
rect 9068 38560 9122 38940
rect 9196 38560 9250 38940
rect 9324 38560 9378 38940
rect 9452 38560 9506 38940
rect 9580 38560 9634 38940
rect 9708 38560 9762 38940
rect 9836 38560 9890 38940
rect 9964 38560 10018 38940
rect 10092 38560 10146 38940
rect 10220 38560 10274 38940
rect 10348 38560 10402 38940
rect 10476 38560 10530 38940
rect 10604 38560 10658 38940
rect 10732 38560 10786 38940
rect 10860 38560 10914 38940
rect 10988 38560 11042 38940
rect 11216 38556 11270 38944
rect 11344 38556 11398 38944
rect 11472 38556 11526 38944
rect 5030 38334 11624 38340
rect 5030 38286 5036 38334
rect 5036 38286 11618 38334
rect 11618 38286 11624 38334
rect 5030 38280 11624 38286
rect 30824 3490 31922 3858
rect 30824 798 31922 1166
<< metal2 >>
rect 5040 39142 5108 39152
rect 11070 39146 11136 39152
rect 5040 39086 5046 39142
rect 5102 39086 5108 39142
rect 5518 39140 5584 39146
rect 5040 39076 5108 39086
rect 5256 39086 5524 39140
rect 5578 39086 5584 39140
rect 11070 39092 11076 39146
rect 11130 39092 11398 39146
rect 11070 39086 11136 39092
rect 5124 38936 5180 38946
rect 5124 38546 5180 38556
rect 5256 38944 5310 39086
rect 5518 39080 5584 39086
rect 5256 38550 5310 38556
rect 5386 38936 5442 38946
rect 5386 38546 5442 38556
rect 5612 38940 5668 38950
rect 5612 38550 5668 38560
rect 5740 38940 5796 38950
rect 5740 38550 5796 38560
rect 5868 38940 5924 38950
rect 5868 38550 5924 38560
rect 5996 38940 6052 38950
rect 5996 38550 6052 38560
rect 6124 38940 6180 38950
rect 6124 38550 6180 38560
rect 6252 38940 6308 38950
rect 6252 38550 6308 38560
rect 6380 38940 6436 38950
rect 6380 38550 6436 38560
rect 6508 38940 6564 38950
rect 6508 38550 6564 38560
rect 6636 38940 6692 38950
rect 6636 38550 6692 38560
rect 6764 38940 6820 38950
rect 6764 38550 6820 38560
rect 6892 38940 6948 38950
rect 6892 38550 6948 38560
rect 7020 38940 7076 38950
rect 7020 38550 7076 38560
rect 7148 38940 7204 38950
rect 7148 38550 7204 38560
rect 7276 38940 7332 38950
rect 7276 38550 7332 38560
rect 7404 38940 7460 38950
rect 7404 38550 7460 38560
rect 7532 38940 7588 38950
rect 7532 38550 7588 38560
rect 7660 38940 7716 38950
rect 7660 38550 7716 38560
rect 7788 38940 7844 38950
rect 7788 38550 7844 38560
rect 7916 38940 7972 38950
rect 7916 38550 7972 38560
rect 8172 38940 8228 38950
rect 8172 38550 8228 38560
rect 8300 38940 8356 38950
rect 8300 38550 8356 38560
rect 8428 38940 8484 38950
rect 8428 38550 8484 38560
rect 8556 38940 8612 38950
rect 8556 38550 8612 38560
rect 8684 38940 8740 38950
rect 8684 38550 8740 38560
rect 8812 38940 8868 38950
rect 8812 38550 8868 38560
rect 8940 38940 8996 38950
rect 8940 38550 8996 38560
rect 9068 38940 9124 38950
rect 9068 38550 9124 38560
rect 9196 38940 9252 38950
rect 9196 38550 9252 38560
rect 9324 38940 9380 38950
rect 9324 38550 9380 38560
rect 9452 38940 9508 38950
rect 9452 38550 9508 38560
rect 9580 38940 9636 38950
rect 9580 38550 9636 38560
rect 9708 38940 9764 38950
rect 9708 38550 9764 38560
rect 9836 38940 9892 38950
rect 9836 38550 9892 38560
rect 9964 38940 10020 38950
rect 9964 38550 10020 38560
rect 10092 38940 10148 38950
rect 10092 38550 10148 38560
rect 10220 38940 10276 38950
rect 10220 38550 10276 38560
rect 10348 38940 10404 38950
rect 10348 38550 10404 38560
rect 10476 38940 10532 38950
rect 10476 38550 10532 38560
rect 10604 38940 10660 38950
rect 10604 38550 10660 38560
rect 10732 38940 10788 38950
rect 10732 38550 10788 38560
rect 10860 38940 10916 38950
rect 10860 38550 10916 38560
rect 10988 38940 11044 38950
rect 10988 38550 11044 38560
rect 11216 38944 11270 38950
rect 11216 38496 11270 38556
rect 11344 38944 11398 39092
rect 11544 39142 11612 39152
rect 11544 39086 11550 39142
rect 11606 39086 11612 39142
rect 11544 39076 11612 39086
rect 11344 38550 11398 38556
rect 11472 38944 11526 38950
rect 11472 38496 11526 38556
rect 11216 38442 31428 38496
rect 11736 38388 31428 38442
rect 5024 38340 11630 38344
rect 5024 38280 5030 38340
rect 11624 38280 11630 38340
rect 5024 38276 11630 38280
rect 31316 3878 31428 38388
rect 30804 3858 31942 3878
rect 30804 3490 30824 3858
rect 31922 3490 31942 3858
rect 30804 3470 31942 3490
rect 30804 1166 31942 1186
rect 30804 798 30824 1166
rect 31922 798 31942 1166
rect 30804 778 31942 798
<< via2 >>
rect 5046 39140 5102 39142
rect 5046 39086 5102 39140
rect 5124 38556 5178 38936
rect 5178 38556 5180 38936
rect 5386 38556 5440 38936
rect 5440 38556 5442 38936
rect 5612 38560 5666 38940
rect 5666 38560 5668 38940
rect 5740 38560 5794 38940
rect 5794 38560 5796 38940
rect 5868 38560 5922 38940
rect 5922 38560 5924 38940
rect 5996 38560 6050 38940
rect 6050 38560 6052 38940
rect 6124 38560 6178 38940
rect 6178 38560 6180 38940
rect 6252 38560 6306 38940
rect 6306 38560 6308 38940
rect 6380 38560 6434 38940
rect 6434 38560 6436 38940
rect 6508 38560 6562 38940
rect 6562 38560 6564 38940
rect 6636 38560 6690 38940
rect 6690 38560 6692 38940
rect 6764 38560 6818 38940
rect 6818 38560 6820 38940
rect 6892 38560 6946 38940
rect 6946 38560 6948 38940
rect 7020 38560 7074 38940
rect 7074 38560 7076 38940
rect 7148 38560 7202 38940
rect 7202 38560 7204 38940
rect 7276 38560 7330 38940
rect 7330 38560 7332 38940
rect 7404 38560 7458 38940
rect 7458 38560 7460 38940
rect 7532 38560 7586 38940
rect 7586 38560 7588 38940
rect 7660 38560 7714 38940
rect 7714 38560 7716 38940
rect 7788 38560 7842 38940
rect 7842 38560 7844 38940
rect 7916 38560 7970 38940
rect 7970 38560 7972 38940
rect 8172 38560 8226 38940
rect 8226 38560 8228 38940
rect 8300 38560 8354 38940
rect 8354 38560 8356 38940
rect 8428 38560 8482 38940
rect 8482 38560 8484 38940
rect 8556 38560 8610 38940
rect 8610 38560 8612 38940
rect 8684 38560 8738 38940
rect 8738 38560 8740 38940
rect 8812 38560 8866 38940
rect 8866 38560 8868 38940
rect 8940 38560 8994 38940
rect 8994 38560 8996 38940
rect 9068 38560 9122 38940
rect 9122 38560 9124 38940
rect 9196 38560 9250 38940
rect 9250 38560 9252 38940
rect 9324 38560 9378 38940
rect 9378 38560 9380 38940
rect 9452 38560 9506 38940
rect 9506 38560 9508 38940
rect 9580 38560 9634 38940
rect 9634 38560 9636 38940
rect 9708 38560 9762 38940
rect 9762 38560 9764 38940
rect 9836 38560 9890 38940
rect 9890 38560 9892 38940
rect 9964 38560 10018 38940
rect 10018 38560 10020 38940
rect 10092 38560 10146 38940
rect 10146 38560 10148 38940
rect 10220 38560 10274 38940
rect 10274 38560 10276 38940
rect 10348 38560 10402 38940
rect 10402 38560 10404 38940
rect 10476 38560 10530 38940
rect 10530 38560 10532 38940
rect 10604 38560 10658 38940
rect 10658 38560 10660 38940
rect 10732 38560 10786 38940
rect 10786 38560 10788 38940
rect 10860 38560 10914 38940
rect 10914 38560 10916 38940
rect 10988 38560 11042 38940
rect 11042 38560 11044 38940
rect 11550 39140 11606 39142
rect 11550 39086 11606 39140
rect 5034 38282 11620 38338
rect 30824 798 31922 1166
<< metal3 >>
rect 11546 40232 11610 40238
rect 11546 40162 11610 40168
rect 5042 40032 5106 40038
rect 5042 39962 5106 39968
rect 300 39840 2300 39850
rect 300 39060 310 39840
rect 890 39060 1710 39840
rect 2290 39060 2300 39840
rect 5044 39148 5104 39962
rect 11548 39148 11608 40162
rect 5040 39142 5108 39148
rect 5040 39086 5046 39142
rect 5102 39086 5108 39142
rect 5040 39080 5108 39086
rect 11544 39142 11612 39148
rect 11544 39086 11550 39142
rect 11606 39086 11612 39142
rect 11544 39080 11612 39086
rect 300 39050 2300 39060
rect 5118 38936 5186 38946
rect 5118 38556 5120 38936
rect 5184 38556 5186 38936
rect 5118 38546 5186 38556
rect 5380 38936 5448 38946
rect 5380 38556 5382 38936
rect 5446 38556 5448 38936
rect 5380 38546 5448 38556
rect 5606 38940 5674 38950
rect 5606 38560 5608 38940
rect 5672 38560 5674 38940
rect 5606 38550 5674 38560
rect 5734 38940 5802 38950
rect 5734 38560 5736 38940
rect 5800 38560 5802 38940
rect 5734 38550 5802 38560
rect 5862 38940 5930 38950
rect 5862 38560 5864 38940
rect 5928 38560 5930 38940
rect 5862 38550 5930 38560
rect 5990 38940 6058 38950
rect 5990 38560 5992 38940
rect 6056 38560 6058 38940
rect 5990 38550 6058 38560
rect 6118 38940 6186 38950
rect 6118 38560 6120 38940
rect 6184 38560 6186 38940
rect 6118 38550 6186 38560
rect 6246 38940 6314 38950
rect 6246 38560 6248 38940
rect 6312 38560 6314 38940
rect 6246 38550 6314 38560
rect 6374 38940 6442 38950
rect 6374 38560 6376 38940
rect 6440 38560 6442 38940
rect 6374 38550 6442 38560
rect 6502 38940 6570 38950
rect 6502 38560 6504 38940
rect 6568 38560 6570 38940
rect 6502 38550 6570 38560
rect 6630 38940 6698 38950
rect 6630 38560 6632 38940
rect 6696 38560 6698 38940
rect 6630 38550 6698 38560
rect 6758 38940 6826 38950
rect 6758 38560 6760 38940
rect 6824 38560 6826 38940
rect 6758 38550 6826 38560
rect 6886 38940 6954 38950
rect 6886 38560 6888 38940
rect 6952 38560 6954 38940
rect 6886 38550 6954 38560
rect 7014 38940 7082 38950
rect 7014 38560 7016 38940
rect 7080 38560 7082 38940
rect 7014 38550 7082 38560
rect 7142 38940 7210 38950
rect 7142 38560 7144 38940
rect 7208 38560 7210 38940
rect 7142 38550 7210 38560
rect 7270 38940 7338 38950
rect 7270 38560 7272 38940
rect 7336 38560 7338 38940
rect 7270 38550 7338 38560
rect 7398 38940 7466 38950
rect 7398 38560 7400 38940
rect 7464 38560 7466 38940
rect 7398 38550 7466 38560
rect 7526 38940 7594 38950
rect 7526 38560 7528 38940
rect 7592 38560 7594 38940
rect 7526 38550 7594 38560
rect 7654 38940 7722 38950
rect 7654 38560 7656 38940
rect 7720 38560 7722 38940
rect 7654 38550 7722 38560
rect 7782 38940 7850 38950
rect 7782 38560 7784 38940
rect 7848 38560 7850 38940
rect 7782 38550 7850 38560
rect 7910 38940 7978 38950
rect 7910 38560 7912 38940
rect 7976 38560 7978 38940
rect 7910 38550 7978 38560
rect 8166 38940 8234 38950
rect 8166 38560 8168 38940
rect 8232 38560 8234 38940
rect 8166 38550 8234 38560
rect 8294 38940 8362 38950
rect 8294 38560 8296 38940
rect 8360 38560 8362 38940
rect 8294 38550 8362 38560
rect 8422 38940 8490 38950
rect 8422 38560 8424 38940
rect 8488 38560 8490 38940
rect 8422 38550 8490 38560
rect 8550 38940 8618 38950
rect 8550 38560 8552 38940
rect 8616 38560 8618 38940
rect 8550 38550 8618 38560
rect 8678 38940 8746 38950
rect 8678 38560 8680 38940
rect 8744 38560 8746 38940
rect 8678 38550 8746 38560
rect 8806 38940 8874 38950
rect 8806 38560 8808 38940
rect 8872 38560 8874 38940
rect 8806 38550 8874 38560
rect 8934 38940 9002 38950
rect 8934 38560 8936 38940
rect 9000 38560 9002 38940
rect 8934 38550 9002 38560
rect 9062 38940 9130 38950
rect 9062 38560 9064 38940
rect 9128 38560 9130 38940
rect 9062 38550 9130 38560
rect 9190 38940 9258 38950
rect 9190 38560 9192 38940
rect 9256 38560 9258 38940
rect 9190 38550 9258 38560
rect 9318 38940 9386 38950
rect 9318 38560 9320 38940
rect 9384 38560 9386 38940
rect 9318 38550 9386 38560
rect 9446 38940 9514 38950
rect 9446 38560 9448 38940
rect 9512 38560 9514 38940
rect 9446 38550 9514 38560
rect 9574 38940 9642 38950
rect 9574 38560 9576 38940
rect 9640 38560 9642 38940
rect 9574 38550 9642 38560
rect 9702 38940 9770 38950
rect 9702 38560 9704 38940
rect 9768 38560 9770 38940
rect 9702 38550 9770 38560
rect 9830 38940 9898 38950
rect 9830 38560 9832 38940
rect 9896 38560 9898 38940
rect 9830 38550 9898 38560
rect 9958 38940 10026 38950
rect 9958 38560 9960 38940
rect 10024 38560 10026 38940
rect 9958 38550 10026 38560
rect 10086 38940 10154 38950
rect 10086 38560 10088 38940
rect 10152 38560 10154 38940
rect 10086 38550 10154 38560
rect 10214 38940 10282 38950
rect 10214 38560 10216 38940
rect 10280 38560 10282 38940
rect 10214 38550 10282 38560
rect 10342 38940 10410 38950
rect 10342 38560 10344 38940
rect 10408 38560 10410 38940
rect 10342 38550 10410 38560
rect 10470 38940 10538 38950
rect 10470 38560 10472 38940
rect 10536 38560 10538 38940
rect 10470 38550 10538 38560
rect 10598 38940 10666 38950
rect 10598 38560 10600 38940
rect 10664 38560 10666 38940
rect 10598 38550 10666 38560
rect 10726 38940 10794 38950
rect 10726 38560 10728 38940
rect 10792 38560 10794 38940
rect 10726 38550 10794 38560
rect 10854 38940 10922 38950
rect 10854 38560 10856 38940
rect 10920 38560 10922 38940
rect 10854 38550 10922 38560
rect 10982 38940 11050 38950
rect 10982 38560 10984 38940
rect 11048 38560 11050 38940
rect 10982 38550 11050 38560
rect 5024 38342 11630 38344
rect 5024 38278 5034 38342
rect 11040 38338 11630 38342
rect 11620 38282 11630 38338
rect 11040 38278 11630 38282
rect 5024 38276 11630 38278
rect 30804 1166 31942 1186
rect 30804 798 30824 1166
rect 31922 798 31942 1166
rect 30804 778 31942 798
<< via3 >>
rect 11546 40168 11610 40232
rect 5042 39968 5106 40032
rect 310 39060 890 39840
rect 1710 39060 2290 39840
rect 5120 38556 5124 38936
rect 5124 38556 5180 38936
rect 5180 38556 5184 38936
rect 5382 38556 5386 38936
rect 5386 38556 5442 38936
rect 5442 38556 5446 38936
rect 5608 38560 5612 38940
rect 5612 38560 5668 38940
rect 5668 38560 5672 38940
rect 5736 38560 5740 38940
rect 5740 38560 5796 38940
rect 5796 38560 5800 38940
rect 5864 38560 5868 38940
rect 5868 38560 5924 38940
rect 5924 38560 5928 38940
rect 5992 38560 5996 38940
rect 5996 38560 6052 38940
rect 6052 38560 6056 38940
rect 6120 38560 6124 38940
rect 6124 38560 6180 38940
rect 6180 38560 6184 38940
rect 6248 38560 6252 38940
rect 6252 38560 6308 38940
rect 6308 38560 6312 38940
rect 6376 38560 6380 38940
rect 6380 38560 6436 38940
rect 6436 38560 6440 38940
rect 6504 38560 6508 38940
rect 6508 38560 6564 38940
rect 6564 38560 6568 38940
rect 6632 38560 6636 38940
rect 6636 38560 6692 38940
rect 6692 38560 6696 38940
rect 6760 38560 6764 38940
rect 6764 38560 6820 38940
rect 6820 38560 6824 38940
rect 6888 38560 6892 38940
rect 6892 38560 6948 38940
rect 6948 38560 6952 38940
rect 7016 38560 7020 38940
rect 7020 38560 7076 38940
rect 7076 38560 7080 38940
rect 7144 38560 7148 38940
rect 7148 38560 7204 38940
rect 7204 38560 7208 38940
rect 7272 38560 7276 38940
rect 7276 38560 7332 38940
rect 7332 38560 7336 38940
rect 7400 38560 7404 38940
rect 7404 38560 7460 38940
rect 7460 38560 7464 38940
rect 7528 38560 7532 38940
rect 7532 38560 7588 38940
rect 7588 38560 7592 38940
rect 7656 38560 7660 38940
rect 7660 38560 7716 38940
rect 7716 38560 7720 38940
rect 7784 38560 7788 38940
rect 7788 38560 7844 38940
rect 7844 38560 7848 38940
rect 7912 38560 7916 38940
rect 7916 38560 7972 38940
rect 7972 38560 7976 38940
rect 8168 38560 8172 38940
rect 8172 38560 8228 38940
rect 8228 38560 8232 38940
rect 8296 38560 8300 38940
rect 8300 38560 8356 38940
rect 8356 38560 8360 38940
rect 8424 38560 8428 38940
rect 8428 38560 8484 38940
rect 8484 38560 8488 38940
rect 8552 38560 8556 38940
rect 8556 38560 8612 38940
rect 8612 38560 8616 38940
rect 8680 38560 8684 38940
rect 8684 38560 8740 38940
rect 8740 38560 8744 38940
rect 8808 38560 8812 38940
rect 8812 38560 8868 38940
rect 8868 38560 8872 38940
rect 8936 38560 8940 38940
rect 8940 38560 8996 38940
rect 8996 38560 9000 38940
rect 9064 38560 9068 38940
rect 9068 38560 9124 38940
rect 9124 38560 9128 38940
rect 9192 38560 9196 38940
rect 9196 38560 9252 38940
rect 9252 38560 9256 38940
rect 9320 38560 9324 38940
rect 9324 38560 9380 38940
rect 9380 38560 9384 38940
rect 9448 38560 9452 38940
rect 9452 38560 9508 38940
rect 9508 38560 9512 38940
rect 9576 38560 9580 38940
rect 9580 38560 9636 38940
rect 9636 38560 9640 38940
rect 9704 38560 9708 38940
rect 9708 38560 9764 38940
rect 9764 38560 9768 38940
rect 9832 38560 9836 38940
rect 9836 38560 9892 38940
rect 9892 38560 9896 38940
rect 9960 38560 9964 38940
rect 9964 38560 10020 38940
rect 10020 38560 10024 38940
rect 10088 38560 10092 38940
rect 10092 38560 10148 38940
rect 10148 38560 10152 38940
rect 10216 38560 10220 38940
rect 10220 38560 10276 38940
rect 10276 38560 10280 38940
rect 10344 38560 10348 38940
rect 10348 38560 10404 38940
rect 10404 38560 10408 38940
rect 10472 38560 10476 38940
rect 10476 38560 10532 38940
rect 10532 38560 10536 38940
rect 10600 38560 10604 38940
rect 10604 38560 10660 38940
rect 10660 38560 10664 38940
rect 10728 38560 10732 38940
rect 10732 38560 10788 38940
rect 10788 38560 10792 38940
rect 10856 38560 10860 38940
rect 10860 38560 10916 38940
rect 10916 38560 10920 38940
rect 10984 38560 10988 38940
rect 10988 38560 11044 38940
rect 11044 38560 11048 38940
rect 5034 38338 11040 38342
rect 5034 38282 11040 38338
rect 5034 38278 11040 38282
rect 30824 798 31922 1166
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 798 44892 17786 44952
rect 1000 44152 1060 44892
rect 300 39840 900 44152
rect 300 39060 310 39840
rect 890 39060 900 39840
rect 300 820 900 39060
rect 1000 38450 1600 44152
rect 11544 40232 11612 40234
rect 11544 40168 11546 40232
rect 11610 40230 11612 40232
rect 22878 40230 22938 45152
rect 11610 40170 22938 40230
rect 11610 40168 11612 40170
rect 11544 40166 11612 40168
rect 5040 40032 5108 40034
rect 5040 39968 5042 40032
rect 5106 40030 5108 40032
rect 23614 40030 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 5106 39970 23674 40030
rect 5106 39968 5108 39970
rect 5040 39966 5108 39968
rect 1700 39840 10922 39850
rect 1700 39060 1710 39840
rect 2290 39060 10922 39840
rect 1700 39050 10922 39060
rect 5118 38936 5186 38946
rect 5118 38556 5120 38936
rect 5184 38556 5186 38936
rect 5118 38450 5186 38556
rect 5380 38936 5448 38946
rect 5380 38556 5382 38936
rect 5446 38556 5448 38936
rect 5380 38450 5448 38556
rect 5606 38940 5674 38950
rect 5606 38560 5608 38940
rect 5672 38560 5674 38940
rect 5606 38450 5674 38560
rect 5734 38940 5802 39050
rect 5734 38560 5736 38940
rect 5800 38560 5802 38940
rect 5734 38550 5802 38560
rect 5862 38940 5930 38950
rect 5862 38560 5864 38940
rect 5928 38560 5930 38940
rect 5862 38450 5930 38560
rect 5990 38940 6058 39050
rect 5990 38560 5992 38940
rect 6056 38560 6058 38940
rect 5990 38550 6058 38560
rect 6118 38940 6186 38950
rect 6118 38560 6120 38940
rect 6184 38560 6186 38940
rect 6118 38450 6186 38560
rect 6246 38940 6314 39050
rect 6246 38560 6248 38940
rect 6312 38560 6314 38940
rect 6246 38550 6314 38560
rect 6374 38940 6442 38950
rect 6374 38560 6376 38940
rect 6440 38560 6442 38940
rect 6374 38450 6442 38560
rect 6502 38940 6570 39050
rect 6502 38560 6504 38940
rect 6568 38560 6570 38940
rect 6502 38550 6570 38560
rect 6630 38940 6698 38950
rect 6630 38560 6632 38940
rect 6696 38560 6698 38940
rect 6630 38450 6698 38560
rect 6758 38940 6826 39050
rect 6758 38560 6760 38940
rect 6824 38560 6826 38940
rect 6758 38550 6826 38560
rect 6886 38940 6954 38950
rect 6886 38560 6888 38940
rect 6952 38560 6954 38940
rect 6886 38450 6954 38560
rect 7014 38940 7082 39050
rect 7014 38560 7016 38940
rect 7080 38560 7082 38940
rect 7014 38550 7082 38560
rect 7142 38940 7210 38950
rect 7142 38560 7144 38940
rect 7208 38560 7210 38940
rect 7142 38450 7210 38560
rect 7270 38940 7338 39050
rect 7270 38560 7272 38940
rect 7336 38560 7338 38940
rect 7270 38550 7338 38560
rect 7398 38940 7466 38950
rect 7398 38560 7400 38940
rect 7464 38560 7466 38940
rect 7398 38450 7466 38560
rect 7526 38940 7594 39050
rect 7526 38560 7528 38940
rect 7592 38560 7594 38940
rect 7526 38550 7594 38560
rect 7654 38940 7722 38950
rect 7654 38560 7656 38940
rect 7720 38560 7722 38940
rect 7654 38450 7722 38560
rect 7782 38940 7850 39050
rect 7782 38560 7784 38940
rect 7848 38560 7850 38940
rect 7782 38550 7850 38560
rect 7910 38940 7978 38950
rect 7910 38560 7912 38940
rect 7976 38560 7978 38940
rect 7910 38450 7978 38560
rect 8166 38940 8234 38950
rect 8166 38560 8168 38940
rect 8232 38560 8234 38940
rect 8166 38450 8234 38560
rect 8294 38940 8362 39050
rect 8294 38560 8296 38940
rect 8360 38560 8362 38940
rect 8294 38550 8362 38560
rect 8422 38940 8490 38950
rect 8422 38560 8424 38940
rect 8488 38560 8490 38940
rect 8422 38450 8490 38560
rect 8550 38940 8618 39050
rect 8550 38560 8552 38940
rect 8616 38560 8618 38940
rect 8550 38550 8618 38560
rect 8678 38940 8746 38950
rect 8678 38560 8680 38940
rect 8744 38560 8746 38940
rect 8678 38450 8746 38560
rect 8806 38940 8874 39050
rect 8806 38560 8808 38940
rect 8872 38560 8874 38940
rect 8806 38550 8874 38560
rect 8934 38940 9002 38950
rect 8934 38560 8936 38940
rect 9000 38560 9002 38940
rect 8934 38450 9002 38560
rect 9062 38940 9130 39050
rect 9062 38560 9064 38940
rect 9128 38560 9130 38940
rect 9062 38550 9130 38560
rect 9190 38940 9258 38950
rect 9190 38560 9192 38940
rect 9256 38560 9258 38940
rect 9190 38450 9258 38560
rect 9318 38940 9386 39050
rect 9318 38560 9320 38940
rect 9384 38560 9386 38940
rect 9318 38550 9386 38560
rect 9446 38940 9514 38950
rect 9446 38560 9448 38940
rect 9512 38560 9514 38940
rect 9446 38450 9514 38560
rect 9574 38940 9642 39050
rect 9574 38560 9576 38940
rect 9640 38560 9642 38940
rect 9574 38550 9642 38560
rect 9702 38940 9770 38950
rect 9702 38560 9704 38940
rect 9768 38560 9770 38940
rect 9702 38450 9770 38560
rect 9830 38940 9898 39050
rect 9830 38560 9832 38940
rect 9896 38560 9898 38940
rect 9830 38550 9898 38560
rect 9958 38940 10026 38950
rect 9958 38560 9960 38940
rect 10024 38560 10026 38940
rect 9958 38450 10026 38560
rect 10086 38940 10154 39050
rect 10086 38560 10088 38940
rect 10152 38560 10154 38940
rect 10086 38550 10154 38560
rect 10214 38940 10282 38950
rect 10214 38560 10216 38940
rect 10280 38560 10282 38940
rect 10214 38450 10282 38560
rect 10342 38940 10410 39050
rect 10342 38560 10344 38940
rect 10408 38560 10410 38940
rect 10342 38550 10410 38560
rect 10470 38940 10538 38950
rect 10470 38560 10472 38940
rect 10536 38560 10538 38940
rect 10470 38450 10538 38560
rect 10598 38940 10666 39050
rect 10598 38560 10600 38940
rect 10664 38560 10666 38940
rect 10598 38550 10666 38560
rect 10726 38940 10794 38950
rect 10726 38560 10728 38940
rect 10792 38560 10794 38940
rect 10726 38450 10794 38560
rect 10854 38940 10922 39050
rect 10854 38560 10856 38940
rect 10920 38560 10922 38940
rect 10854 38550 10922 38560
rect 10982 38940 11050 38950
rect 10982 38560 10984 38940
rect 11048 38560 11050 38940
rect 10982 38450 11050 38560
rect 1000 38342 11050 38450
rect 1000 38278 5034 38342
rect 11040 38278 11050 38342
rect 1000 37650 11050 38278
rect 1000 1180 1600 37650
rect 1000 1000 27046 1180
rect 300 640 22630 820
rect 9204 200 18214 380
rect 400 0 520 200
rect 4816 0 4936 200
rect 9204 0 9384 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 640
rect 26866 0 27046 1000
rect 30804 1166 31942 1186
rect 30804 798 30824 1166
rect 31922 798 31942 1166
rect 30804 778 31942 798
rect 31282 0 31462 778
use sky130_fd_pr__nfet_01v8_HH22ET  sky130_fd_pr__nfet_01v8_HH22ET_0
timestamp 1713626126
transform 1 0 8327 0 1 38750
box -2855 -410 2855 410
use sky130_fd_pr__nfet_01v8_HX7DH9  sky130_fd_pr__nfet_01v8_HX7DH9_0
timestamp 1713626233
transform 1 0 11371 0 1 38750
box -295 -410 295 410
use sky130_fd_pr__nfet_01v8_HX7DH9  sky130_fd_pr__nfet_01v8_HX7DH9_1
timestamp 1713626233
transform 1 0 5283 0 1 38750
box -295 -410 295 410
use sky130_fd_pr__res_high_po_5p73_VFSSNU  sky130_fd_pr__res_high_po_5p73_VFSSNU_0
timestamp 1713626469
transform 1 0 31373 0 1 2328
box -739 -1728 739 1728
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 600 1000 900 44152 1 FreeSans 720 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 1000 1000 1300 44152 1 FreeSans 720 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
