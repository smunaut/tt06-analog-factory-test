magic
tech sky130A
magscale 1 2
timestamp 1713626126
<< error_p >>
rect -2655 272 -2593 278
rect -2527 272 -2465 278
rect -2399 272 -2337 278
rect -2271 272 -2209 278
rect -2143 272 -2081 278
rect -2015 272 -1953 278
rect -1887 272 -1825 278
rect -1759 272 -1697 278
rect -1631 272 -1569 278
rect -1503 272 -1441 278
rect -1375 272 -1313 278
rect -1247 272 -1185 278
rect -1119 272 -1057 278
rect -991 272 -929 278
rect -863 272 -801 278
rect -735 272 -673 278
rect -607 272 -545 278
rect -479 272 -417 278
rect -351 272 -289 278
rect -223 272 -161 278
rect -95 272 -33 278
rect 33 272 95 278
rect 161 272 223 278
rect 289 272 351 278
rect 417 272 479 278
rect 545 272 607 278
rect 673 272 735 278
rect 801 272 863 278
rect 929 272 991 278
rect 1057 272 1119 278
rect 1185 272 1247 278
rect 1313 272 1375 278
rect 1441 272 1503 278
rect 1569 272 1631 278
rect 1697 272 1759 278
rect 1825 272 1887 278
rect 1953 272 2015 278
rect 2081 272 2143 278
rect 2209 272 2271 278
rect 2337 272 2399 278
rect 2465 272 2527 278
rect 2593 272 2655 278
rect -2655 238 -2643 272
rect -2527 238 -2515 272
rect -2399 238 -2387 272
rect -2271 238 -2259 272
rect -2143 238 -2131 272
rect -2015 238 -2003 272
rect -1887 238 -1875 272
rect -1759 238 -1747 272
rect -1631 238 -1619 272
rect -1503 238 -1491 272
rect -1375 238 -1363 272
rect -1247 238 -1235 272
rect -1119 238 -1107 272
rect -991 238 -979 272
rect -863 238 -851 272
rect -735 238 -723 272
rect -607 238 -595 272
rect -479 238 -467 272
rect -351 238 -339 272
rect -223 238 -211 272
rect -95 238 -83 272
rect 33 238 45 272
rect 161 238 173 272
rect 289 238 301 272
rect 417 238 429 272
rect 545 238 557 272
rect 673 238 685 272
rect 801 238 813 272
rect 929 238 941 272
rect 1057 238 1069 272
rect 1185 238 1197 272
rect 1313 238 1325 272
rect 1441 238 1453 272
rect 1569 238 1581 272
rect 1697 238 1709 272
rect 1825 238 1837 272
rect 1953 238 1965 272
rect 2081 238 2093 272
rect 2209 238 2221 272
rect 2337 238 2349 272
rect 2465 238 2477 272
rect 2593 238 2605 272
rect -2655 232 -2593 238
rect -2527 232 -2465 238
rect -2399 232 -2337 238
rect -2271 232 -2209 238
rect -2143 232 -2081 238
rect -2015 232 -1953 238
rect -1887 232 -1825 238
rect -1759 232 -1697 238
rect -1631 232 -1569 238
rect -1503 232 -1441 238
rect -1375 232 -1313 238
rect -1247 232 -1185 238
rect -1119 232 -1057 238
rect -991 232 -929 238
rect -863 232 -801 238
rect -735 232 -673 238
rect -607 232 -545 238
rect -479 232 -417 238
rect -351 232 -289 238
rect -223 232 -161 238
rect -95 232 -33 238
rect 33 232 95 238
rect 161 232 223 238
rect 289 232 351 238
rect 417 232 479 238
rect 545 232 607 238
rect 673 232 735 238
rect 801 232 863 238
rect 929 232 991 238
rect 1057 232 1119 238
rect 1185 232 1247 238
rect 1313 232 1375 238
rect 1441 232 1503 238
rect 1569 232 1631 238
rect 1697 232 1759 238
rect 1825 232 1887 238
rect 1953 232 2015 238
rect 2081 232 2143 238
rect 2209 232 2271 238
rect 2337 232 2399 238
rect 2465 232 2527 238
rect 2593 232 2655 238
rect -2655 -238 -2593 -232
rect -2527 -238 -2465 -232
rect -2399 -238 -2337 -232
rect -2271 -238 -2209 -232
rect -2143 -238 -2081 -232
rect -2015 -238 -1953 -232
rect -1887 -238 -1825 -232
rect -1759 -238 -1697 -232
rect -1631 -238 -1569 -232
rect -1503 -238 -1441 -232
rect -1375 -238 -1313 -232
rect -1247 -238 -1185 -232
rect -1119 -238 -1057 -232
rect -991 -238 -929 -232
rect -863 -238 -801 -232
rect -735 -238 -673 -232
rect -607 -238 -545 -232
rect -479 -238 -417 -232
rect -351 -238 -289 -232
rect -223 -238 -161 -232
rect -95 -238 -33 -232
rect 33 -238 95 -232
rect 161 -238 223 -232
rect 289 -238 351 -232
rect 417 -238 479 -232
rect 545 -238 607 -232
rect 673 -238 735 -232
rect 801 -238 863 -232
rect 929 -238 991 -232
rect 1057 -238 1119 -232
rect 1185 -238 1247 -232
rect 1313 -238 1375 -232
rect 1441 -238 1503 -232
rect 1569 -238 1631 -232
rect 1697 -238 1759 -232
rect 1825 -238 1887 -232
rect 1953 -238 2015 -232
rect 2081 -238 2143 -232
rect 2209 -238 2271 -232
rect 2337 -238 2399 -232
rect 2465 -238 2527 -232
rect 2593 -238 2655 -232
rect -2655 -272 -2643 -238
rect -2527 -272 -2515 -238
rect -2399 -272 -2387 -238
rect -2271 -272 -2259 -238
rect -2143 -272 -2131 -238
rect -2015 -272 -2003 -238
rect -1887 -272 -1875 -238
rect -1759 -272 -1747 -238
rect -1631 -272 -1619 -238
rect -1503 -272 -1491 -238
rect -1375 -272 -1363 -238
rect -1247 -272 -1235 -238
rect -1119 -272 -1107 -238
rect -991 -272 -979 -238
rect -863 -272 -851 -238
rect -735 -272 -723 -238
rect -607 -272 -595 -238
rect -479 -272 -467 -238
rect -351 -272 -339 -238
rect -223 -272 -211 -238
rect -95 -272 -83 -238
rect 33 -272 45 -238
rect 161 -272 173 -238
rect 289 -272 301 -238
rect 417 -272 429 -238
rect 545 -272 557 -238
rect 673 -272 685 -238
rect 801 -272 813 -238
rect 929 -272 941 -238
rect 1057 -272 1069 -238
rect 1185 -272 1197 -238
rect 1313 -272 1325 -238
rect 1441 -272 1453 -238
rect 1569 -272 1581 -238
rect 1697 -272 1709 -238
rect 1825 -272 1837 -238
rect 1953 -272 1965 -238
rect 2081 -272 2093 -238
rect 2209 -272 2221 -238
rect 2337 -272 2349 -238
rect 2465 -272 2477 -238
rect 2593 -272 2605 -238
rect -2655 -278 -2593 -272
rect -2527 -278 -2465 -272
rect -2399 -278 -2337 -272
rect -2271 -278 -2209 -272
rect -2143 -278 -2081 -272
rect -2015 -278 -1953 -272
rect -1887 -278 -1825 -272
rect -1759 -278 -1697 -272
rect -1631 -278 -1569 -272
rect -1503 -278 -1441 -272
rect -1375 -278 -1313 -272
rect -1247 -278 -1185 -272
rect -1119 -278 -1057 -272
rect -991 -278 -929 -272
rect -863 -278 -801 -272
rect -735 -278 -673 -272
rect -607 -278 -545 -272
rect -479 -278 -417 -272
rect -351 -278 -289 -272
rect -223 -278 -161 -272
rect -95 -278 -33 -272
rect 33 -278 95 -272
rect 161 -278 223 -272
rect 289 -278 351 -272
rect 417 -278 479 -272
rect 545 -278 607 -272
rect 673 -278 735 -272
rect 801 -278 863 -272
rect 929 -278 991 -272
rect 1057 -278 1119 -272
rect 1185 -278 1247 -272
rect 1313 -278 1375 -272
rect 1441 -278 1503 -272
rect 1569 -278 1631 -272
rect 1697 -278 1759 -272
rect 1825 -278 1887 -272
rect 1953 -278 2015 -272
rect 2081 -278 2143 -272
rect 2209 -278 2271 -272
rect 2337 -278 2399 -272
rect 2465 -278 2527 -272
rect 2593 -278 2655 -272
<< pwell >>
rect -2855 -410 2855 410
<< nmos >>
rect -2659 -200 -2589 200
rect -2531 -200 -2461 200
rect -2403 -200 -2333 200
rect -2275 -200 -2205 200
rect -2147 -200 -2077 200
rect -2019 -200 -1949 200
rect -1891 -200 -1821 200
rect -1763 -200 -1693 200
rect -1635 -200 -1565 200
rect -1507 -200 -1437 200
rect -1379 -200 -1309 200
rect -1251 -200 -1181 200
rect -1123 -200 -1053 200
rect -995 -200 -925 200
rect -867 -200 -797 200
rect -739 -200 -669 200
rect -611 -200 -541 200
rect -483 -200 -413 200
rect -355 -200 -285 200
rect -227 -200 -157 200
rect -99 -200 -29 200
rect 29 -200 99 200
rect 157 -200 227 200
rect 285 -200 355 200
rect 413 -200 483 200
rect 541 -200 611 200
rect 669 -200 739 200
rect 797 -200 867 200
rect 925 -200 995 200
rect 1053 -200 1123 200
rect 1181 -200 1251 200
rect 1309 -200 1379 200
rect 1437 -200 1507 200
rect 1565 -200 1635 200
rect 1693 -200 1763 200
rect 1821 -200 1891 200
rect 1949 -200 2019 200
rect 2077 -200 2147 200
rect 2205 -200 2275 200
rect 2333 -200 2403 200
rect 2461 -200 2531 200
rect 2589 -200 2659 200
<< ndiff >>
rect -2717 188 -2659 200
rect -2717 -188 -2705 188
rect -2671 -188 -2659 188
rect -2717 -200 -2659 -188
rect -2589 188 -2531 200
rect -2589 -188 -2577 188
rect -2543 -188 -2531 188
rect -2589 -200 -2531 -188
rect -2461 188 -2403 200
rect -2461 -188 -2449 188
rect -2415 -188 -2403 188
rect -2461 -200 -2403 -188
rect -2333 188 -2275 200
rect -2333 -188 -2321 188
rect -2287 -188 -2275 188
rect -2333 -200 -2275 -188
rect -2205 188 -2147 200
rect -2205 -188 -2193 188
rect -2159 -188 -2147 188
rect -2205 -200 -2147 -188
rect -2077 188 -2019 200
rect -2077 -188 -2065 188
rect -2031 -188 -2019 188
rect -2077 -200 -2019 -188
rect -1949 188 -1891 200
rect -1949 -188 -1937 188
rect -1903 -188 -1891 188
rect -1949 -200 -1891 -188
rect -1821 188 -1763 200
rect -1821 -188 -1809 188
rect -1775 -188 -1763 188
rect -1821 -200 -1763 -188
rect -1693 188 -1635 200
rect -1693 -188 -1681 188
rect -1647 -188 -1635 188
rect -1693 -200 -1635 -188
rect -1565 188 -1507 200
rect -1565 -188 -1553 188
rect -1519 -188 -1507 188
rect -1565 -200 -1507 -188
rect -1437 188 -1379 200
rect -1437 -188 -1425 188
rect -1391 -188 -1379 188
rect -1437 -200 -1379 -188
rect -1309 188 -1251 200
rect -1309 -188 -1297 188
rect -1263 -188 -1251 188
rect -1309 -200 -1251 -188
rect -1181 188 -1123 200
rect -1181 -188 -1169 188
rect -1135 -188 -1123 188
rect -1181 -200 -1123 -188
rect -1053 188 -995 200
rect -1053 -188 -1041 188
rect -1007 -188 -995 188
rect -1053 -200 -995 -188
rect -925 188 -867 200
rect -925 -188 -913 188
rect -879 -188 -867 188
rect -925 -200 -867 -188
rect -797 188 -739 200
rect -797 -188 -785 188
rect -751 -188 -739 188
rect -797 -200 -739 -188
rect -669 188 -611 200
rect -669 -188 -657 188
rect -623 -188 -611 188
rect -669 -200 -611 -188
rect -541 188 -483 200
rect -541 -188 -529 188
rect -495 -188 -483 188
rect -541 -200 -483 -188
rect -413 188 -355 200
rect -413 -188 -401 188
rect -367 -188 -355 188
rect -413 -200 -355 -188
rect -285 188 -227 200
rect -285 -188 -273 188
rect -239 -188 -227 188
rect -285 -200 -227 -188
rect -157 188 -99 200
rect -157 -188 -145 188
rect -111 -188 -99 188
rect -157 -200 -99 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 99 188 157 200
rect 99 -188 111 188
rect 145 -188 157 188
rect 99 -200 157 -188
rect 227 188 285 200
rect 227 -188 239 188
rect 273 -188 285 188
rect 227 -200 285 -188
rect 355 188 413 200
rect 355 -188 367 188
rect 401 -188 413 188
rect 355 -200 413 -188
rect 483 188 541 200
rect 483 -188 495 188
rect 529 -188 541 188
rect 483 -200 541 -188
rect 611 188 669 200
rect 611 -188 623 188
rect 657 -188 669 188
rect 611 -200 669 -188
rect 739 188 797 200
rect 739 -188 751 188
rect 785 -188 797 188
rect 739 -200 797 -188
rect 867 188 925 200
rect 867 -188 879 188
rect 913 -188 925 188
rect 867 -200 925 -188
rect 995 188 1053 200
rect 995 -188 1007 188
rect 1041 -188 1053 188
rect 995 -200 1053 -188
rect 1123 188 1181 200
rect 1123 -188 1135 188
rect 1169 -188 1181 188
rect 1123 -200 1181 -188
rect 1251 188 1309 200
rect 1251 -188 1263 188
rect 1297 -188 1309 188
rect 1251 -200 1309 -188
rect 1379 188 1437 200
rect 1379 -188 1391 188
rect 1425 -188 1437 188
rect 1379 -200 1437 -188
rect 1507 188 1565 200
rect 1507 -188 1519 188
rect 1553 -188 1565 188
rect 1507 -200 1565 -188
rect 1635 188 1693 200
rect 1635 -188 1647 188
rect 1681 -188 1693 188
rect 1635 -200 1693 -188
rect 1763 188 1821 200
rect 1763 -188 1775 188
rect 1809 -188 1821 188
rect 1763 -200 1821 -188
rect 1891 188 1949 200
rect 1891 -188 1903 188
rect 1937 -188 1949 188
rect 1891 -200 1949 -188
rect 2019 188 2077 200
rect 2019 -188 2031 188
rect 2065 -188 2077 188
rect 2019 -200 2077 -188
rect 2147 188 2205 200
rect 2147 -188 2159 188
rect 2193 -188 2205 188
rect 2147 -200 2205 -188
rect 2275 188 2333 200
rect 2275 -188 2287 188
rect 2321 -188 2333 188
rect 2275 -200 2333 -188
rect 2403 188 2461 200
rect 2403 -188 2415 188
rect 2449 -188 2461 188
rect 2403 -200 2461 -188
rect 2531 188 2589 200
rect 2531 -188 2543 188
rect 2577 -188 2589 188
rect 2531 -200 2589 -188
rect 2659 188 2717 200
rect 2659 -188 2671 188
rect 2705 -188 2717 188
rect 2659 -200 2717 -188
<< ndiffc >>
rect -2705 -188 -2671 188
rect -2577 -188 -2543 188
rect -2449 -188 -2415 188
rect -2321 -188 -2287 188
rect -2193 -188 -2159 188
rect -2065 -188 -2031 188
rect -1937 -188 -1903 188
rect -1809 -188 -1775 188
rect -1681 -188 -1647 188
rect -1553 -188 -1519 188
rect -1425 -188 -1391 188
rect -1297 -188 -1263 188
rect -1169 -188 -1135 188
rect -1041 -188 -1007 188
rect -913 -188 -879 188
rect -785 -188 -751 188
rect -657 -188 -623 188
rect -529 -188 -495 188
rect -401 -188 -367 188
rect -273 -188 -239 188
rect -145 -188 -111 188
rect -17 -188 17 188
rect 111 -188 145 188
rect 239 -188 273 188
rect 367 -188 401 188
rect 495 -188 529 188
rect 623 -188 657 188
rect 751 -188 785 188
rect 879 -188 913 188
rect 1007 -188 1041 188
rect 1135 -188 1169 188
rect 1263 -188 1297 188
rect 1391 -188 1425 188
rect 1519 -188 1553 188
rect 1647 -188 1681 188
rect 1775 -188 1809 188
rect 1903 -188 1937 188
rect 2031 -188 2065 188
rect 2159 -188 2193 188
rect 2287 -188 2321 188
rect 2415 -188 2449 188
rect 2543 -188 2577 188
rect 2671 -188 2705 188
<< psubdiff >>
rect -2819 340 -2723 374
rect 2723 340 2819 374
rect -2819 278 -2785 340
rect 2785 278 2819 340
rect -2819 -340 -2785 -278
rect 2785 -340 2819 -278
rect -2819 -374 -2723 -340
rect 2723 -374 2819 -340
<< psubdiffcont >>
rect -2723 340 2723 374
rect -2819 -278 -2785 278
rect 2785 -278 2819 278
rect -2723 -374 2723 -340
<< poly >>
rect -2659 272 -2589 288
rect -2659 238 -2643 272
rect -2605 238 -2589 272
rect -2659 200 -2589 238
rect -2531 272 -2461 288
rect -2531 238 -2515 272
rect -2477 238 -2461 272
rect -2531 200 -2461 238
rect -2403 272 -2333 288
rect -2403 238 -2387 272
rect -2349 238 -2333 272
rect -2403 200 -2333 238
rect -2275 272 -2205 288
rect -2275 238 -2259 272
rect -2221 238 -2205 272
rect -2275 200 -2205 238
rect -2147 272 -2077 288
rect -2147 238 -2131 272
rect -2093 238 -2077 272
rect -2147 200 -2077 238
rect -2019 272 -1949 288
rect -2019 238 -2003 272
rect -1965 238 -1949 272
rect -2019 200 -1949 238
rect -1891 272 -1821 288
rect -1891 238 -1875 272
rect -1837 238 -1821 272
rect -1891 200 -1821 238
rect -1763 272 -1693 288
rect -1763 238 -1747 272
rect -1709 238 -1693 272
rect -1763 200 -1693 238
rect -1635 272 -1565 288
rect -1635 238 -1619 272
rect -1581 238 -1565 272
rect -1635 200 -1565 238
rect -1507 272 -1437 288
rect -1507 238 -1491 272
rect -1453 238 -1437 272
rect -1507 200 -1437 238
rect -1379 272 -1309 288
rect -1379 238 -1363 272
rect -1325 238 -1309 272
rect -1379 200 -1309 238
rect -1251 272 -1181 288
rect -1251 238 -1235 272
rect -1197 238 -1181 272
rect -1251 200 -1181 238
rect -1123 272 -1053 288
rect -1123 238 -1107 272
rect -1069 238 -1053 272
rect -1123 200 -1053 238
rect -995 272 -925 288
rect -995 238 -979 272
rect -941 238 -925 272
rect -995 200 -925 238
rect -867 272 -797 288
rect -867 238 -851 272
rect -813 238 -797 272
rect -867 200 -797 238
rect -739 272 -669 288
rect -739 238 -723 272
rect -685 238 -669 272
rect -739 200 -669 238
rect -611 272 -541 288
rect -611 238 -595 272
rect -557 238 -541 272
rect -611 200 -541 238
rect -483 272 -413 288
rect -483 238 -467 272
rect -429 238 -413 272
rect -483 200 -413 238
rect -355 272 -285 288
rect -355 238 -339 272
rect -301 238 -285 272
rect -355 200 -285 238
rect -227 272 -157 288
rect -227 238 -211 272
rect -173 238 -157 272
rect -227 200 -157 238
rect -99 272 -29 288
rect -99 238 -83 272
rect -45 238 -29 272
rect -99 200 -29 238
rect 29 272 99 288
rect 29 238 45 272
rect 83 238 99 272
rect 29 200 99 238
rect 157 272 227 288
rect 157 238 173 272
rect 211 238 227 272
rect 157 200 227 238
rect 285 272 355 288
rect 285 238 301 272
rect 339 238 355 272
rect 285 200 355 238
rect 413 272 483 288
rect 413 238 429 272
rect 467 238 483 272
rect 413 200 483 238
rect 541 272 611 288
rect 541 238 557 272
rect 595 238 611 272
rect 541 200 611 238
rect 669 272 739 288
rect 669 238 685 272
rect 723 238 739 272
rect 669 200 739 238
rect 797 272 867 288
rect 797 238 813 272
rect 851 238 867 272
rect 797 200 867 238
rect 925 272 995 288
rect 925 238 941 272
rect 979 238 995 272
rect 925 200 995 238
rect 1053 272 1123 288
rect 1053 238 1069 272
rect 1107 238 1123 272
rect 1053 200 1123 238
rect 1181 272 1251 288
rect 1181 238 1197 272
rect 1235 238 1251 272
rect 1181 200 1251 238
rect 1309 272 1379 288
rect 1309 238 1325 272
rect 1363 238 1379 272
rect 1309 200 1379 238
rect 1437 272 1507 288
rect 1437 238 1453 272
rect 1491 238 1507 272
rect 1437 200 1507 238
rect 1565 272 1635 288
rect 1565 238 1581 272
rect 1619 238 1635 272
rect 1565 200 1635 238
rect 1693 272 1763 288
rect 1693 238 1709 272
rect 1747 238 1763 272
rect 1693 200 1763 238
rect 1821 272 1891 288
rect 1821 238 1837 272
rect 1875 238 1891 272
rect 1821 200 1891 238
rect 1949 272 2019 288
rect 1949 238 1965 272
rect 2003 238 2019 272
rect 1949 200 2019 238
rect 2077 272 2147 288
rect 2077 238 2093 272
rect 2131 238 2147 272
rect 2077 200 2147 238
rect 2205 272 2275 288
rect 2205 238 2221 272
rect 2259 238 2275 272
rect 2205 200 2275 238
rect 2333 272 2403 288
rect 2333 238 2349 272
rect 2387 238 2403 272
rect 2333 200 2403 238
rect 2461 272 2531 288
rect 2461 238 2477 272
rect 2515 238 2531 272
rect 2461 200 2531 238
rect 2589 272 2659 288
rect 2589 238 2605 272
rect 2643 238 2659 272
rect 2589 200 2659 238
rect -2659 -238 -2589 -200
rect -2659 -272 -2643 -238
rect -2605 -272 -2589 -238
rect -2659 -288 -2589 -272
rect -2531 -238 -2461 -200
rect -2531 -272 -2515 -238
rect -2477 -272 -2461 -238
rect -2531 -288 -2461 -272
rect -2403 -238 -2333 -200
rect -2403 -272 -2387 -238
rect -2349 -272 -2333 -238
rect -2403 -288 -2333 -272
rect -2275 -238 -2205 -200
rect -2275 -272 -2259 -238
rect -2221 -272 -2205 -238
rect -2275 -288 -2205 -272
rect -2147 -238 -2077 -200
rect -2147 -272 -2131 -238
rect -2093 -272 -2077 -238
rect -2147 -288 -2077 -272
rect -2019 -238 -1949 -200
rect -2019 -272 -2003 -238
rect -1965 -272 -1949 -238
rect -2019 -288 -1949 -272
rect -1891 -238 -1821 -200
rect -1891 -272 -1875 -238
rect -1837 -272 -1821 -238
rect -1891 -288 -1821 -272
rect -1763 -238 -1693 -200
rect -1763 -272 -1747 -238
rect -1709 -272 -1693 -238
rect -1763 -288 -1693 -272
rect -1635 -238 -1565 -200
rect -1635 -272 -1619 -238
rect -1581 -272 -1565 -238
rect -1635 -288 -1565 -272
rect -1507 -238 -1437 -200
rect -1507 -272 -1491 -238
rect -1453 -272 -1437 -238
rect -1507 -288 -1437 -272
rect -1379 -238 -1309 -200
rect -1379 -272 -1363 -238
rect -1325 -272 -1309 -238
rect -1379 -288 -1309 -272
rect -1251 -238 -1181 -200
rect -1251 -272 -1235 -238
rect -1197 -272 -1181 -238
rect -1251 -288 -1181 -272
rect -1123 -238 -1053 -200
rect -1123 -272 -1107 -238
rect -1069 -272 -1053 -238
rect -1123 -288 -1053 -272
rect -995 -238 -925 -200
rect -995 -272 -979 -238
rect -941 -272 -925 -238
rect -995 -288 -925 -272
rect -867 -238 -797 -200
rect -867 -272 -851 -238
rect -813 -272 -797 -238
rect -867 -288 -797 -272
rect -739 -238 -669 -200
rect -739 -272 -723 -238
rect -685 -272 -669 -238
rect -739 -288 -669 -272
rect -611 -238 -541 -200
rect -611 -272 -595 -238
rect -557 -272 -541 -238
rect -611 -288 -541 -272
rect -483 -238 -413 -200
rect -483 -272 -467 -238
rect -429 -272 -413 -238
rect -483 -288 -413 -272
rect -355 -238 -285 -200
rect -355 -272 -339 -238
rect -301 -272 -285 -238
rect -355 -288 -285 -272
rect -227 -238 -157 -200
rect -227 -272 -211 -238
rect -173 -272 -157 -238
rect -227 -288 -157 -272
rect -99 -238 -29 -200
rect -99 -272 -83 -238
rect -45 -272 -29 -238
rect -99 -288 -29 -272
rect 29 -238 99 -200
rect 29 -272 45 -238
rect 83 -272 99 -238
rect 29 -288 99 -272
rect 157 -238 227 -200
rect 157 -272 173 -238
rect 211 -272 227 -238
rect 157 -288 227 -272
rect 285 -238 355 -200
rect 285 -272 301 -238
rect 339 -272 355 -238
rect 285 -288 355 -272
rect 413 -238 483 -200
rect 413 -272 429 -238
rect 467 -272 483 -238
rect 413 -288 483 -272
rect 541 -238 611 -200
rect 541 -272 557 -238
rect 595 -272 611 -238
rect 541 -288 611 -272
rect 669 -238 739 -200
rect 669 -272 685 -238
rect 723 -272 739 -238
rect 669 -288 739 -272
rect 797 -238 867 -200
rect 797 -272 813 -238
rect 851 -272 867 -238
rect 797 -288 867 -272
rect 925 -238 995 -200
rect 925 -272 941 -238
rect 979 -272 995 -238
rect 925 -288 995 -272
rect 1053 -238 1123 -200
rect 1053 -272 1069 -238
rect 1107 -272 1123 -238
rect 1053 -288 1123 -272
rect 1181 -238 1251 -200
rect 1181 -272 1197 -238
rect 1235 -272 1251 -238
rect 1181 -288 1251 -272
rect 1309 -238 1379 -200
rect 1309 -272 1325 -238
rect 1363 -272 1379 -238
rect 1309 -288 1379 -272
rect 1437 -238 1507 -200
rect 1437 -272 1453 -238
rect 1491 -272 1507 -238
rect 1437 -288 1507 -272
rect 1565 -238 1635 -200
rect 1565 -272 1581 -238
rect 1619 -272 1635 -238
rect 1565 -288 1635 -272
rect 1693 -238 1763 -200
rect 1693 -272 1709 -238
rect 1747 -272 1763 -238
rect 1693 -288 1763 -272
rect 1821 -238 1891 -200
rect 1821 -272 1837 -238
rect 1875 -272 1891 -238
rect 1821 -288 1891 -272
rect 1949 -238 2019 -200
rect 1949 -272 1965 -238
rect 2003 -272 2019 -238
rect 1949 -288 2019 -272
rect 2077 -238 2147 -200
rect 2077 -272 2093 -238
rect 2131 -272 2147 -238
rect 2077 -288 2147 -272
rect 2205 -238 2275 -200
rect 2205 -272 2221 -238
rect 2259 -272 2275 -238
rect 2205 -288 2275 -272
rect 2333 -238 2403 -200
rect 2333 -272 2349 -238
rect 2387 -272 2403 -238
rect 2333 -288 2403 -272
rect 2461 -238 2531 -200
rect 2461 -272 2477 -238
rect 2515 -272 2531 -238
rect 2461 -288 2531 -272
rect 2589 -238 2659 -200
rect 2589 -272 2605 -238
rect 2643 -272 2659 -238
rect 2589 -288 2659 -272
<< polycont >>
rect -2643 238 -2605 272
rect -2515 238 -2477 272
rect -2387 238 -2349 272
rect -2259 238 -2221 272
rect -2131 238 -2093 272
rect -2003 238 -1965 272
rect -1875 238 -1837 272
rect -1747 238 -1709 272
rect -1619 238 -1581 272
rect -1491 238 -1453 272
rect -1363 238 -1325 272
rect -1235 238 -1197 272
rect -1107 238 -1069 272
rect -979 238 -941 272
rect -851 238 -813 272
rect -723 238 -685 272
rect -595 238 -557 272
rect -467 238 -429 272
rect -339 238 -301 272
rect -211 238 -173 272
rect -83 238 -45 272
rect 45 238 83 272
rect 173 238 211 272
rect 301 238 339 272
rect 429 238 467 272
rect 557 238 595 272
rect 685 238 723 272
rect 813 238 851 272
rect 941 238 979 272
rect 1069 238 1107 272
rect 1197 238 1235 272
rect 1325 238 1363 272
rect 1453 238 1491 272
rect 1581 238 1619 272
rect 1709 238 1747 272
rect 1837 238 1875 272
rect 1965 238 2003 272
rect 2093 238 2131 272
rect 2221 238 2259 272
rect 2349 238 2387 272
rect 2477 238 2515 272
rect 2605 238 2643 272
rect -2643 -272 -2605 -238
rect -2515 -272 -2477 -238
rect -2387 -272 -2349 -238
rect -2259 -272 -2221 -238
rect -2131 -272 -2093 -238
rect -2003 -272 -1965 -238
rect -1875 -272 -1837 -238
rect -1747 -272 -1709 -238
rect -1619 -272 -1581 -238
rect -1491 -272 -1453 -238
rect -1363 -272 -1325 -238
rect -1235 -272 -1197 -238
rect -1107 -272 -1069 -238
rect -979 -272 -941 -238
rect -851 -272 -813 -238
rect -723 -272 -685 -238
rect -595 -272 -557 -238
rect -467 -272 -429 -238
rect -339 -272 -301 -238
rect -211 -272 -173 -238
rect -83 -272 -45 -238
rect 45 -272 83 -238
rect 173 -272 211 -238
rect 301 -272 339 -238
rect 429 -272 467 -238
rect 557 -272 595 -238
rect 685 -272 723 -238
rect 813 -272 851 -238
rect 941 -272 979 -238
rect 1069 -272 1107 -238
rect 1197 -272 1235 -238
rect 1325 -272 1363 -238
rect 1453 -272 1491 -238
rect 1581 -272 1619 -238
rect 1709 -272 1747 -238
rect 1837 -272 1875 -238
rect 1965 -272 2003 -238
rect 2093 -272 2131 -238
rect 2221 -272 2259 -238
rect 2349 -272 2387 -238
rect 2477 -272 2515 -238
rect 2605 -272 2643 -238
<< locali >>
rect -2819 340 -2723 374
rect 2723 340 2819 374
rect -2819 278 -2785 340
rect 2785 278 2819 340
rect -2659 238 -2643 272
rect -2605 238 -2589 272
rect -2531 238 -2515 272
rect -2477 238 -2461 272
rect -2403 238 -2387 272
rect -2349 238 -2333 272
rect -2275 238 -2259 272
rect -2221 238 -2205 272
rect -2147 238 -2131 272
rect -2093 238 -2077 272
rect -2019 238 -2003 272
rect -1965 238 -1949 272
rect -1891 238 -1875 272
rect -1837 238 -1821 272
rect -1763 238 -1747 272
rect -1709 238 -1693 272
rect -1635 238 -1619 272
rect -1581 238 -1565 272
rect -1507 238 -1491 272
rect -1453 238 -1437 272
rect -1379 238 -1363 272
rect -1325 238 -1309 272
rect -1251 238 -1235 272
rect -1197 238 -1181 272
rect -1123 238 -1107 272
rect -1069 238 -1053 272
rect -995 238 -979 272
rect -941 238 -925 272
rect -867 238 -851 272
rect -813 238 -797 272
rect -739 238 -723 272
rect -685 238 -669 272
rect -611 238 -595 272
rect -557 238 -541 272
rect -483 238 -467 272
rect -429 238 -413 272
rect -355 238 -339 272
rect -301 238 -285 272
rect -227 238 -211 272
rect -173 238 -157 272
rect -99 238 -83 272
rect -45 238 -29 272
rect 29 238 45 272
rect 83 238 99 272
rect 157 238 173 272
rect 211 238 227 272
rect 285 238 301 272
rect 339 238 355 272
rect 413 238 429 272
rect 467 238 483 272
rect 541 238 557 272
rect 595 238 611 272
rect 669 238 685 272
rect 723 238 739 272
rect 797 238 813 272
rect 851 238 867 272
rect 925 238 941 272
rect 979 238 995 272
rect 1053 238 1069 272
rect 1107 238 1123 272
rect 1181 238 1197 272
rect 1235 238 1251 272
rect 1309 238 1325 272
rect 1363 238 1379 272
rect 1437 238 1453 272
rect 1491 238 1507 272
rect 1565 238 1581 272
rect 1619 238 1635 272
rect 1693 238 1709 272
rect 1747 238 1763 272
rect 1821 238 1837 272
rect 1875 238 1891 272
rect 1949 238 1965 272
rect 2003 238 2019 272
rect 2077 238 2093 272
rect 2131 238 2147 272
rect 2205 238 2221 272
rect 2259 238 2275 272
rect 2333 238 2349 272
rect 2387 238 2403 272
rect 2461 238 2477 272
rect 2515 238 2531 272
rect 2589 238 2605 272
rect 2643 238 2659 272
rect -2705 188 -2671 204
rect -2705 -204 -2671 -188
rect -2577 188 -2543 204
rect -2577 -204 -2543 -188
rect -2449 188 -2415 204
rect -2449 -204 -2415 -188
rect -2321 188 -2287 204
rect -2321 -204 -2287 -188
rect -2193 188 -2159 204
rect -2193 -204 -2159 -188
rect -2065 188 -2031 204
rect -2065 -204 -2031 -188
rect -1937 188 -1903 204
rect -1937 -204 -1903 -188
rect -1809 188 -1775 204
rect -1809 -204 -1775 -188
rect -1681 188 -1647 204
rect -1681 -204 -1647 -188
rect -1553 188 -1519 204
rect -1553 -204 -1519 -188
rect -1425 188 -1391 204
rect -1425 -204 -1391 -188
rect -1297 188 -1263 204
rect -1297 -204 -1263 -188
rect -1169 188 -1135 204
rect -1169 -204 -1135 -188
rect -1041 188 -1007 204
rect -1041 -204 -1007 -188
rect -913 188 -879 204
rect -913 -204 -879 -188
rect -785 188 -751 204
rect -785 -204 -751 -188
rect -657 188 -623 204
rect -657 -204 -623 -188
rect -529 188 -495 204
rect -529 -204 -495 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -273 188 -239 204
rect -273 -204 -239 -188
rect -145 188 -111 204
rect -145 -204 -111 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 111 188 145 204
rect 111 -204 145 -188
rect 239 188 273 204
rect 239 -204 273 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 495 188 529 204
rect 495 -204 529 -188
rect 623 188 657 204
rect 623 -204 657 -188
rect 751 188 785 204
rect 751 -204 785 -188
rect 879 188 913 204
rect 879 -204 913 -188
rect 1007 188 1041 204
rect 1007 -204 1041 -188
rect 1135 188 1169 204
rect 1135 -204 1169 -188
rect 1263 188 1297 204
rect 1263 -204 1297 -188
rect 1391 188 1425 204
rect 1391 -204 1425 -188
rect 1519 188 1553 204
rect 1519 -204 1553 -188
rect 1647 188 1681 204
rect 1647 -204 1681 -188
rect 1775 188 1809 204
rect 1775 -204 1809 -188
rect 1903 188 1937 204
rect 1903 -204 1937 -188
rect 2031 188 2065 204
rect 2031 -204 2065 -188
rect 2159 188 2193 204
rect 2159 -204 2193 -188
rect 2287 188 2321 204
rect 2287 -204 2321 -188
rect 2415 188 2449 204
rect 2415 -204 2449 -188
rect 2543 188 2577 204
rect 2543 -204 2577 -188
rect 2671 188 2705 204
rect 2671 -204 2705 -188
rect -2659 -272 -2643 -238
rect -2605 -272 -2589 -238
rect -2531 -272 -2515 -238
rect -2477 -272 -2461 -238
rect -2403 -272 -2387 -238
rect -2349 -272 -2333 -238
rect -2275 -272 -2259 -238
rect -2221 -272 -2205 -238
rect -2147 -272 -2131 -238
rect -2093 -272 -2077 -238
rect -2019 -272 -2003 -238
rect -1965 -272 -1949 -238
rect -1891 -272 -1875 -238
rect -1837 -272 -1821 -238
rect -1763 -272 -1747 -238
rect -1709 -272 -1693 -238
rect -1635 -272 -1619 -238
rect -1581 -272 -1565 -238
rect -1507 -272 -1491 -238
rect -1453 -272 -1437 -238
rect -1379 -272 -1363 -238
rect -1325 -272 -1309 -238
rect -1251 -272 -1235 -238
rect -1197 -272 -1181 -238
rect -1123 -272 -1107 -238
rect -1069 -272 -1053 -238
rect -995 -272 -979 -238
rect -941 -272 -925 -238
rect -867 -272 -851 -238
rect -813 -272 -797 -238
rect -739 -272 -723 -238
rect -685 -272 -669 -238
rect -611 -272 -595 -238
rect -557 -272 -541 -238
rect -483 -272 -467 -238
rect -429 -272 -413 -238
rect -355 -272 -339 -238
rect -301 -272 -285 -238
rect -227 -272 -211 -238
rect -173 -272 -157 -238
rect -99 -272 -83 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 83 -272 99 -238
rect 157 -272 173 -238
rect 211 -272 227 -238
rect 285 -272 301 -238
rect 339 -272 355 -238
rect 413 -272 429 -238
rect 467 -272 483 -238
rect 541 -272 557 -238
rect 595 -272 611 -238
rect 669 -272 685 -238
rect 723 -272 739 -238
rect 797 -272 813 -238
rect 851 -272 867 -238
rect 925 -272 941 -238
rect 979 -272 995 -238
rect 1053 -272 1069 -238
rect 1107 -272 1123 -238
rect 1181 -272 1197 -238
rect 1235 -272 1251 -238
rect 1309 -272 1325 -238
rect 1363 -272 1379 -238
rect 1437 -272 1453 -238
rect 1491 -272 1507 -238
rect 1565 -272 1581 -238
rect 1619 -272 1635 -238
rect 1693 -272 1709 -238
rect 1747 -272 1763 -238
rect 1821 -272 1837 -238
rect 1875 -272 1891 -238
rect 1949 -272 1965 -238
rect 2003 -272 2019 -238
rect 2077 -272 2093 -238
rect 2131 -272 2147 -238
rect 2205 -272 2221 -238
rect 2259 -272 2275 -238
rect 2333 -272 2349 -238
rect 2387 -272 2403 -238
rect 2461 -272 2477 -238
rect 2515 -272 2531 -238
rect 2589 -272 2605 -238
rect 2643 -272 2659 -238
rect -2819 -340 -2785 -278
rect 2785 -340 2819 -278
rect -2819 -374 -2723 -340
rect 2723 -374 2819 -340
<< viali >>
rect -2643 238 -2605 272
rect -2515 238 -2477 272
rect -2387 238 -2349 272
rect -2259 238 -2221 272
rect -2131 238 -2093 272
rect -2003 238 -1965 272
rect -1875 238 -1837 272
rect -1747 238 -1709 272
rect -1619 238 -1581 272
rect -1491 238 -1453 272
rect -1363 238 -1325 272
rect -1235 238 -1197 272
rect -1107 238 -1069 272
rect -979 238 -941 272
rect -851 238 -813 272
rect -723 238 -685 272
rect -595 238 -557 272
rect -467 238 -429 272
rect -339 238 -301 272
rect -211 238 -173 272
rect -83 238 -45 272
rect 45 238 83 272
rect 173 238 211 272
rect 301 238 339 272
rect 429 238 467 272
rect 557 238 595 272
rect 685 238 723 272
rect 813 238 851 272
rect 941 238 979 272
rect 1069 238 1107 272
rect 1197 238 1235 272
rect 1325 238 1363 272
rect 1453 238 1491 272
rect 1581 238 1619 272
rect 1709 238 1747 272
rect 1837 238 1875 272
rect 1965 238 2003 272
rect 2093 238 2131 272
rect 2221 238 2259 272
rect 2349 238 2387 272
rect 2477 238 2515 272
rect 2605 238 2643 272
rect -2705 -188 -2671 188
rect -2577 -188 -2543 188
rect -2449 -188 -2415 188
rect -2321 -188 -2287 188
rect -2193 -188 -2159 188
rect -2065 -188 -2031 188
rect -1937 -188 -1903 188
rect -1809 -188 -1775 188
rect -1681 -188 -1647 188
rect -1553 -188 -1519 188
rect -1425 -188 -1391 188
rect -1297 -188 -1263 188
rect -1169 -188 -1135 188
rect -1041 -188 -1007 188
rect -913 -188 -879 188
rect -785 -188 -751 188
rect -657 -188 -623 188
rect -529 -188 -495 188
rect -401 -188 -367 188
rect -273 -188 -239 188
rect -145 -188 -111 188
rect -17 -188 17 188
rect 111 -188 145 188
rect 239 -188 273 188
rect 367 -188 401 188
rect 495 -188 529 188
rect 623 -188 657 188
rect 751 -188 785 188
rect 879 -188 913 188
rect 1007 -188 1041 188
rect 1135 -188 1169 188
rect 1263 -188 1297 188
rect 1391 -188 1425 188
rect 1519 -188 1553 188
rect 1647 -188 1681 188
rect 1775 -188 1809 188
rect 1903 -188 1937 188
rect 2031 -188 2065 188
rect 2159 -188 2193 188
rect 2287 -188 2321 188
rect 2415 -188 2449 188
rect 2543 -188 2577 188
rect 2671 -188 2705 188
rect -2643 -272 -2605 -238
rect -2515 -272 -2477 -238
rect -2387 -272 -2349 -238
rect -2259 -272 -2221 -238
rect -2131 -272 -2093 -238
rect -2003 -272 -1965 -238
rect -1875 -272 -1837 -238
rect -1747 -272 -1709 -238
rect -1619 -272 -1581 -238
rect -1491 -272 -1453 -238
rect -1363 -272 -1325 -238
rect -1235 -272 -1197 -238
rect -1107 -272 -1069 -238
rect -979 -272 -941 -238
rect -851 -272 -813 -238
rect -723 -272 -685 -238
rect -595 -272 -557 -238
rect -467 -272 -429 -238
rect -339 -272 -301 -238
rect -211 -272 -173 -238
rect -83 -272 -45 -238
rect 45 -272 83 -238
rect 173 -272 211 -238
rect 301 -272 339 -238
rect 429 -272 467 -238
rect 557 -272 595 -238
rect 685 -272 723 -238
rect 813 -272 851 -238
rect 941 -272 979 -238
rect 1069 -272 1107 -238
rect 1197 -272 1235 -238
rect 1325 -272 1363 -238
rect 1453 -272 1491 -238
rect 1581 -272 1619 -238
rect 1709 -272 1747 -238
rect 1837 -272 1875 -238
rect 1965 -272 2003 -238
rect 2093 -272 2131 -238
rect 2221 -272 2259 -238
rect 2349 -272 2387 -238
rect 2477 -272 2515 -238
rect 2605 -272 2643 -238
<< metal1 >>
rect -2655 272 -2593 278
rect -2655 238 -2643 272
rect -2605 238 -2593 272
rect -2655 232 -2593 238
rect -2527 272 -2465 278
rect -2527 238 -2515 272
rect -2477 238 -2465 272
rect -2527 232 -2465 238
rect -2399 272 -2337 278
rect -2399 238 -2387 272
rect -2349 238 -2337 272
rect -2399 232 -2337 238
rect -2271 272 -2209 278
rect -2271 238 -2259 272
rect -2221 238 -2209 272
rect -2271 232 -2209 238
rect -2143 272 -2081 278
rect -2143 238 -2131 272
rect -2093 238 -2081 272
rect -2143 232 -2081 238
rect -2015 272 -1953 278
rect -2015 238 -2003 272
rect -1965 238 -1953 272
rect -2015 232 -1953 238
rect -1887 272 -1825 278
rect -1887 238 -1875 272
rect -1837 238 -1825 272
rect -1887 232 -1825 238
rect -1759 272 -1697 278
rect -1759 238 -1747 272
rect -1709 238 -1697 272
rect -1759 232 -1697 238
rect -1631 272 -1569 278
rect -1631 238 -1619 272
rect -1581 238 -1569 272
rect -1631 232 -1569 238
rect -1503 272 -1441 278
rect -1503 238 -1491 272
rect -1453 238 -1441 272
rect -1503 232 -1441 238
rect -1375 272 -1313 278
rect -1375 238 -1363 272
rect -1325 238 -1313 272
rect -1375 232 -1313 238
rect -1247 272 -1185 278
rect -1247 238 -1235 272
rect -1197 238 -1185 272
rect -1247 232 -1185 238
rect -1119 272 -1057 278
rect -1119 238 -1107 272
rect -1069 238 -1057 272
rect -1119 232 -1057 238
rect -991 272 -929 278
rect -991 238 -979 272
rect -941 238 -929 272
rect -991 232 -929 238
rect -863 272 -801 278
rect -863 238 -851 272
rect -813 238 -801 272
rect -863 232 -801 238
rect -735 272 -673 278
rect -735 238 -723 272
rect -685 238 -673 272
rect -735 232 -673 238
rect -607 272 -545 278
rect -607 238 -595 272
rect -557 238 -545 272
rect -607 232 -545 238
rect -479 272 -417 278
rect -479 238 -467 272
rect -429 238 -417 272
rect -479 232 -417 238
rect -351 272 -289 278
rect -351 238 -339 272
rect -301 238 -289 272
rect -351 232 -289 238
rect -223 272 -161 278
rect -223 238 -211 272
rect -173 238 -161 272
rect -223 232 -161 238
rect -95 272 -33 278
rect -95 238 -83 272
rect -45 238 -33 272
rect -95 232 -33 238
rect 33 272 95 278
rect 33 238 45 272
rect 83 238 95 272
rect 33 232 95 238
rect 161 272 223 278
rect 161 238 173 272
rect 211 238 223 272
rect 161 232 223 238
rect 289 272 351 278
rect 289 238 301 272
rect 339 238 351 272
rect 289 232 351 238
rect 417 272 479 278
rect 417 238 429 272
rect 467 238 479 272
rect 417 232 479 238
rect 545 272 607 278
rect 545 238 557 272
rect 595 238 607 272
rect 545 232 607 238
rect 673 272 735 278
rect 673 238 685 272
rect 723 238 735 272
rect 673 232 735 238
rect 801 272 863 278
rect 801 238 813 272
rect 851 238 863 272
rect 801 232 863 238
rect 929 272 991 278
rect 929 238 941 272
rect 979 238 991 272
rect 929 232 991 238
rect 1057 272 1119 278
rect 1057 238 1069 272
rect 1107 238 1119 272
rect 1057 232 1119 238
rect 1185 272 1247 278
rect 1185 238 1197 272
rect 1235 238 1247 272
rect 1185 232 1247 238
rect 1313 272 1375 278
rect 1313 238 1325 272
rect 1363 238 1375 272
rect 1313 232 1375 238
rect 1441 272 1503 278
rect 1441 238 1453 272
rect 1491 238 1503 272
rect 1441 232 1503 238
rect 1569 272 1631 278
rect 1569 238 1581 272
rect 1619 238 1631 272
rect 1569 232 1631 238
rect 1697 272 1759 278
rect 1697 238 1709 272
rect 1747 238 1759 272
rect 1697 232 1759 238
rect 1825 272 1887 278
rect 1825 238 1837 272
rect 1875 238 1887 272
rect 1825 232 1887 238
rect 1953 272 2015 278
rect 1953 238 1965 272
rect 2003 238 2015 272
rect 1953 232 2015 238
rect 2081 272 2143 278
rect 2081 238 2093 272
rect 2131 238 2143 272
rect 2081 232 2143 238
rect 2209 272 2271 278
rect 2209 238 2221 272
rect 2259 238 2271 272
rect 2209 232 2271 238
rect 2337 272 2399 278
rect 2337 238 2349 272
rect 2387 238 2399 272
rect 2337 232 2399 238
rect 2465 272 2527 278
rect 2465 238 2477 272
rect 2515 238 2527 272
rect 2465 232 2527 238
rect 2593 272 2655 278
rect 2593 238 2605 272
rect 2643 238 2655 272
rect 2593 232 2655 238
rect -2711 188 -2665 200
rect -2711 -188 -2705 188
rect -2671 -188 -2665 188
rect -2711 -200 -2665 -188
rect -2583 188 -2537 200
rect -2583 -188 -2577 188
rect -2543 -188 -2537 188
rect -2583 -200 -2537 -188
rect -2455 188 -2409 200
rect -2455 -188 -2449 188
rect -2415 -188 -2409 188
rect -2455 -200 -2409 -188
rect -2327 188 -2281 200
rect -2327 -188 -2321 188
rect -2287 -188 -2281 188
rect -2327 -200 -2281 -188
rect -2199 188 -2153 200
rect -2199 -188 -2193 188
rect -2159 -188 -2153 188
rect -2199 -200 -2153 -188
rect -2071 188 -2025 200
rect -2071 -188 -2065 188
rect -2031 -188 -2025 188
rect -2071 -200 -2025 -188
rect -1943 188 -1897 200
rect -1943 -188 -1937 188
rect -1903 -188 -1897 188
rect -1943 -200 -1897 -188
rect -1815 188 -1769 200
rect -1815 -188 -1809 188
rect -1775 -188 -1769 188
rect -1815 -200 -1769 -188
rect -1687 188 -1641 200
rect -1687 -188 -1681 188
rect -1647 -188 -1641 188
rect -1687 -200 -1641 -188
rect -1559 188 -1513 200
rect -1559 -188 -1553 188
rect -1519 -188 -1513 188
rect -1559 -200 -1513 -188
rect -1431 188 -1385 200
rect -1431 -188 -1425 188
rect -1391 -188 -1385 188
rect -1431 -200 -1385 -188
rect -1303 188 -1257 200
rect -1303 -188 -1297 188
rect -1263 -188 -1257 188
rect -1303 -200 -1257 -188
rect -1175 188 -1129 200
rect -1175 -188 -1169 188
rect -1135 -188 -1129 188
rect -1175 -200 -1129 -188
rect -1047 188 -1001 200
rect -1047 -188 -1041 188
rect -1007 -188 -1001 188
rect -1047 -200 -1001 -188
rect -919 188 -873 200
rect -919 -188 -913 188
rect -879 -188 -873 188
rect -919 -200 -873 -188
rect -791 188 -745 200
rect -791 -188 -785 188
rect -751 -188 -745 188
rect -791 -200 -745 -188
rect -663 188 -617 200
rect -663 -188 -657 188
rect -623 -188 -617 188
rect -663 -200 -617 -188
rect -535 188 -489 200
rect -535 -188 -529 188
rect -495 -188 -489 188
rect -535 -200 -489 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -279 188 -233 200
rect -279 -188 -273 188
rect -239 -188 -233 188
rect -279 -200 -233 -188
rect -151 188 -105 200
rect -151 -188 -145 188
rect -111 -188 -105 188
rect -151 -200 -105 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 105 188 151 200
rect 105 -188 111 188
rect 145 -188 151 188
rect 105 -200 151 -188
rect 233 188 279 200
rect 233 -188 239 188
rect 273 -188 279 188
rect 233 -200 279 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 489 188 535 200
rect 489 -188 495 188
rect 529 -188 535 188
rect 489 -200 535 -188
rect 617 188 663 200
rect 617 -188 623 188
rect 657 -188 663 188
rect 617 -200 663 -188
rect 745 188 791 200
rect 745 -188 751 188
rect 785 -188 791 188
rect 745 -200 791 -188
rect 873 188 919 200
rect 873 -188 879 188
rect 913 -188 919 188
rect 873 -200 919 -188
rect 1001 188 1047 200
rect 1001 -188 1007 188
rect 1041 -188 1047 188
rect 1001 -200 1047 -188
rect 1129 188 1175 200
rect 1129 -188 1135 188
rect 1169 -188 1175 188
rect 1129 -200 1175 -188
rect 1257 188 1303 200
rect 1257 -188 1263 188
rect 1297 -188 1303 188
rect 1257 -200 1303 -188
rect 1385 188 1431 200
rect 1385 -188 1391 188
rect 1425 -188 1431 188
rect 1385 -200 1431 -188
rect 1513 188 1559 200
rect 1513 -188 1519 188
rect 1553 -188 1559 188
rect 1513 -200 1559 -188
rect 1641 188 1687 200
rect 1641 -188 1647 188
rect 1681 -188 1687 188
rect 1641 -200 1687 -188
rect 1769 188 1815 200
rect 1769 -188 1775 188
rect 1809 -188 1815 188
rect 1769 -200 1815 -188
rect 1897 188 1943 200
rect 1897 -188 1903 188
rect 1937 -188 1943 188
rect 1897 -200 1943 -188
rect 2025 188 2071 200
rect 2025 -188 2031 188
rect 2065 -188 2071 188
rect 2025 -200 2071 -188
rect 2153 188 2199 200
rect 2153 -188 2159 188
rect 2193 -188 2199 188
rect 2153 -200 2199 -188
rect 2281 188 2327 200
rect 2281 -188 2287 188
rect 2321 -188 2327 188
rect 2281 -200 2327 -188
rect 2409 188 2455 200
rect 2409 -188 2415 188
rect 2449 -188 2455 188
rect 2409 -200 2455 -188
rect 2537 188 2583 200
rect 2537 -188 2543 188
rect 2577 -188 2583 188
rect 2537 -200 2583 -188
rect 2665 188 2711 200
rect 2665 -188 2671 188
rect 2705 -188 2711 188
rect 2665 -200 2711 -188
rect -2655 -238 -2593 -232
rect -2655 -272 -2643 -238
rect -2605 -272 -2593 -238
rect -2655 -278 -2593 -272
rect -2527 -238 -2465 -232
rect -2527 -272 -2515 -238
rect -2477 -272 -2465 -238
rect -2527 -278 -2465 -272
rect -2399 -238 -2337 -232
rect -2399 -272 -2387 -238
rect -2349 -272 -2337 -238
rect -2399 -278 -2337 -272
rect -2271 -238 -2209 -232
rect -2271 -272 -2259 -238
rect -2221 -272 -2209 -238
rect -2271 -278 -2209 -272
rect -2143 -238 -2081 -232
rect -2143 -272 -2131 -238
rect -2093 -272 -2081 -238
rect -2143 -278 -2081 -272
rect -2015 -238 -1953 -232
rect -2015 -272 -2003 -238
rect -1965 -272 -1953 -238
rect -2015 -278 -1953 -272
rect -1887 -238 -1825 -232
rect -1887 -272 -1875 -238
rect -1837 -272 -1825 -238
rect -1887 -278 -1825 -272
rect -1759 -238 -1697 -232
rect -1759 -272 -1747 -238
rect -1709 -272 -1697 -238
rect -1759 -278 -1697 -272
rect -1631 -238 -1569 -232
rect -1631 -272 -1619 -238
rect -1581 -272 -1569 -238
rect -1631 -278 -1569 -272
rect -1503 -238 -1441 -232
rect -1503 -272 -1491 -238
rect -1453 -272 -1441 -238
rect -1503 -278 -1441 -272
rect -1375 -238 -1313 -232
rect -1375 -272 -1363 -238
rect -1325 -272 -1313 -238
rect -1375 -278 -1313 -272
rect -1247 -238 -1185 -232
rect -1247 -272 -1235 -238
rect -1197 -272 -1185 -238
rect -1247 -278 -1185 -272
rect -1119 -238 -1057 -232
rect -1119 -272 -1107 -238
rect -1069 -272 -1057 -238
rect -1119 -278 -1057 -272
rect -991 -238 -929 -232
rect -991 -272 -979 -238
rect -941 -272 -929 -238
rect -991 -278 -929 -272
rect -863 -238 -801 -232
rect -863 -272 -851 -238
rect -813 -272 -801 -238
rect -863 -278 -801 -272
rect -735 -238 -673 -232
rect -735 -272 -723 -238
rect -685 -272 -673 -238
rect -735 -278 -673 -272
rect -607 -238 -545 -232
rect -607 -272 -595 -238
rect -557 -272 -545 -238
rect -607 -278 -545 -272
rect -479 -238 -417 -232
rect -479 -272 -467 -238
rect -429 -272 -417 -238
rect -479 -278 -417 -272
rect -351 -238 -289 -232
rect -351 -272 -339 -238
rect -301 -272 -289 -238
rect -351 -278 -289 -272
rect -223 -238 -161 -232
rect -223 -272 -211 -238
rect -173 -272 -161 -238
rect -223 -278 -161 -272
rect -95 -238 -33 -232
rect -95 -272 -83 -238
rect -45 -272 -33 -238
rect -95 -278 -33 -272
rect 33 -238 95 -232
rect 33 -272 45 -238
rect 83 -272 95 -238
rect 33 -278 95 -272
rect 161 -238 223 -232
rect 161 -272 173 -238
rect 211 -272 223 -238
rect 161 -278 223 -272
rect 289 -238 351 -232
rect 289 -272 301 -238
rect 339 -272 351 -238
rect 289 -278 351 -272
rect 417 -238 479 -232
rect 417 -272 429 -238
rect 467 -272 479 -238
rect 417 -278 479 -272
rect 545 -238 607 -232
rect 545 -272 557 -238
rect 595 -272 607 -238
rect 545 -278 607 -272
rect 673 -238 735 -232
rect 673 -272 685 -238
rect 723 -272 735 -238
rect 673 -278 735 -272
rect 801 -238 863 -232
rect 801 -272 813 -238
rect 851 -272 863 -238
rect 801 -278 863 -272
rect 929 -238 991 -232
rect 929 -272 941 -238
rect 979 -272 991 -238
rect 929 -278 991 -272
rect 1057 -238 1119 -232
rect 1057 -272 1069 -238
rect 1107 -272 1119 -238
rect 1057 -278 1119 -272
rect 1185 -238 1247 -232
rect 1185 -272 1197 -238
rect 1235 -272 1247 -238
rect 1185 -278 1247 -272
rect 1313 -238 1375 -232
rect 1313 -272 1325 -238
rect 1363 -272 1375 -238
rect 1313 -278 1375 -272
rect 1441 -238 1503 -232
rect 1441 -272 1453 -238
rect 1491 -272 1503 -238
rect 1441 -278 1503 -272
rect 1569 -238 1631 -232
rect 1569 -272 1581 -238
rect 1619 -272 1631 -238
rect 1569 -278 1631 -272
rect 1697 -238 1759 -232
rect 1697 -272 1709 -238
rect 1747 -272 1759 -238
rect 1697 -278 1759 -272
rect 1825 -238 1887 -232
rect 1825 -272 1837 -238
rect 1875 -272 1887 -238
rect 1825 -278 1887 -272
rect 1953 -238 2015 -232
rect 1953 -272 1965 -238
rect 2003 -272 2015 -238
rect 1953 -278 2015 -272
rect 2081 -238 2143 -232
rect 2081 -272 2093 -238
rect 2131 -272 2143 -238
rect 2081 -278 2143 -272
rect 2209 -238 2271 -232
rect 2209 -272 2221 -238
rect 2259 -272 2271 -238
rect 2209 -278 2271 -272
rect 2337 -238 2399 -232
rect 2337 -272 2349 -238
rect 2387 -272 2399 -238
rect 2337 -278 2399 -272
rect 2465 -238 2527 -232
rect 2465 -272 2477 -238
rect 2515 -272 2527 -238
rect 2465 -278 2527 -272
rect 2593 -238 2655 -232
rect 2593 -272 2605 -238
rect 2643 -272 2655 -238
rect 2593 -278 2655 -272
<< properties >>
string FIXED_BBOX -2802 -357 2802 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.35 m 1 nf 42 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
