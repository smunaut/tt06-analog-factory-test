magic
tech sky130A
magscale 1 2
timestamp 1713626233
<< error_p >>
rect -95 272 -33 278
rect 33 272 95 278
rect -95 238 -83 272
rect 33 238 45 272
rect -95 232 -33 238
rect 33 232 95 238
rect -95 -238 -33 -232
rect 33 -238 95 -232
rect -95 -272 -83 -238
rect 33 -272 45 -238
rect -95 -278 -33 -272
rect 33 -278 95 -272
<< pwell >>
rect -295 -410 295 410
<< nmos >>
rect -99 -200 -29 200
rect 29 -200 99 200
<< ndiff >>
rect -157 188 -99 200
rect -157 -188 -145 188
rect -111 -188 -99 188
rect -157 -200 -99 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 99 188 157 200
rect 99 -188 111 188
rect 145 -188 157 188
rect 99 -200 157 -188
<< ndiffc >>
rect -145 -188 -111 188
rect -17 -188 17 188
rect 111 -188 145 188
<< psubdiff >>
rect -259 340 -163 374
rect 163 340 259 374
rect -259 278 -225 340
rect 225 278 259 340
rect -259 -340 -225 -278
rect 225 -340 259 -278
rect -259 -374 -163 -340
rect 163 -374 259 -340
<< psubdiffcont >>
rect -163 340 163 374
rect -259 -278 -225 278
rect 225 -278 259 278
rect -163 -374 163 -340
<< poly >>
rect -99 272 -29 288
rect -99 238 -83 272
rect -45 238 -29 272
rect -99 200 -29 238
rect 29 272 99 288
rect 29 238 45 272
rect 83 238 99 272
rect 29 200 99 238
rect -99 -238 -29 -200
rect -99 -272 -83 -238
rect -45 -272 -29 -238
rect -99 -288 -29 -272
rect 29 -238 99 -200
rect 29 -272 45 -238
rect 83 -272 99 -238
rect 29 -288 99 -272
<< polycont >>
rect -83 238 -45 272
rect 45 238 83 272
rect -83 -272 -45 -238
rect 45 -272 83 -238
<< locali >>
rect -259 340 -163 374
rect 163 340 259 374
rect -259 278 -225 340
rect 225 278 259 340
rect -99 238 -83 272
rect -45 238 -29 272
rect 29 238 45 272
rect 83 238 99 272
rect -145 188 -111 204
rect -145 -204 -111 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 111 188 145 204
rect 111 -204 145 -188
rect -99 -272 -83 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 83 -272 99 -238
rect -259 -340 -225 -278
rect 225 -340 259 -278
rect -259 -374 -163 -340
rect 163 -374 259 -340
<< viali >>
rect -83 238 -45 272
rect 45 238 83 272
rect -145 -188 -111 188
rect -17 -188 17 188
rect 111 -188 145 188
rect -83 -272 -45 -238
rect 45 -272 83 -238
<< metal1 >>
rect -95 272 -33 278
rect -95 238 -83 272
rect -45 238 -33 272
rect -95 232 -33 238
rect 33 272 95 278
rect 33 238 45 272
rect 83 238 95 272
rect 33 232 95 238
rect -151 188 -105 200
rect -151 -188 -145 188
rect -111 -188 -105 188
rect -151 -200 -105 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 105 188 151 200
rect 105 -188 111 188
rect 145 -188 151 188
rect 105 -200 151 -188
rect -95 -238 -33 -232
rect -95 -272 -83 -238
rect -45 -272 -33 -238
rect -95 -278 -33 -272
rect 33 -238 95 -232
rect 33 -272 45 -238
rect 83 -272 95 -238
rect 33 -278 95 -272
<< properties >>
string FIXED_BBOX -242 -357 242 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.35 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
